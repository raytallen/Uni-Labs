module FSM(clk, );

endmodule